/******************************
* file   : bin2bcd.v
* date   : 2019-08-24
* author : lanjunjie250@outlook.com 
******************************/

module bin2bcd(


);



endmodule //bin2bcd