/******************************
* file   : bin2bcd.v
* date   : 2019-08-24
* author : lanjunjie250@outlook.com 
******************************/

module bin2bcd(
    rst_n,
    clk,
    start_en,
    busy_o,

);



endmodule //bin2bcd