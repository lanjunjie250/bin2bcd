/*********************************
* file 	 : top.v
* date   : 2019-08-24
* auther : lanjunjie250@outlook.com
*********************************/

module top();

initial begin
    $display("this is top level");
    $finish;
end

endmodule //top
